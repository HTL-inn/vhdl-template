-- Title: 
-- File: tb_main.vhd
-- Author: 
-- Date: 
-- Description: 

library std;
  use std.textio.all;
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
  --use ieee.std_logic_textio.all; -- not compatible with ghdl
library work;
  use work.main_pkg.all;
  use work.tb_main_pkg.all;
  --use work.std_logic_textio.all; -- not compatible with ghdl
  
-- entity

entity tb_main is
  generic (
    
  );
end tb_main
  
-- architecture `behavior`

architecture behavior of tb_main is
  
begin

end behavior;
