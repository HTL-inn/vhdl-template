-- Title: 
-- File: main_pkg.vhd
-- Author: 
-- Date: 
-- Description: 

library ieee;
  use ieee.std_logic_1164.all;
library work;

-- constants

-- package body

package body main_pkg is
end main_pkg;
