-- Title: 
-- File: main.vhd
-- Author: 
-- Date: 
-- Description: 

library	ieee;
  use ieee.std_logic_1164.all;
library work;

-- entity

entity main is
  generic (
    
  );
  
  port (
      
  );
end main;

-- architecture `behavior`

architecture behavior of main is
  
begin

end behavior
