-- Title: 
-- File: tb_main_pkg.vhd
-- Author: 
-- Date: 
-- Description: 

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
library work;
  use work.DE0_pkg.all;
  use work.main_pkg.all;
  
-- entity

entity tb_main is
  generic (
    
  );
end tb_main;
  
-- architecture `behavior`

architecture behavior of tb_main is
  
begin

end behavior;

-- package

package tb_main_pkg is
  
end tb_main_pkg;

-- package body

package body tb_edge_detector_pkg is
end tb_edge_detector_pkg;
